`include "quadra.vh"


`ifndef LUT_SV
	`define LUT_SV
module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = '0;
        7'b0000001 :  a = '0;
        7'b0000010 :  a = '0;
        7'b0000011 :  a = '0;
        7'b0000100 :  a = '0;
        7'b0000101 :  a = '0;
        7'b0000110 :  a = '0;
        7'b0000111 :  a = '0;
        7'b0001000 :  a = '0;
        7'b0001001 :  a = '0;
        7'b0001010 :  a = '0;
        7'b0001011 :  a = '0;
        7'b0001100 :  a = '0;
        7'b0001101 :  a = '0;
        7'b0001110 :  a = '0;
        7'b0001111 :  a = '0;
        7'b0010000 :  a = '0;
        7'b0010001 :  a = '0;
        7'b0010010 :  a = '0;
        7'b0010011 :  a = '0;
        7'b0010100 :  a = '0;
        7'b0010101 :  a = '0;
        7'b0010110 :  a = '0;
        7'b0010111 :  a = '0;
        7'b0011000 :  a = '0;
        7'b0011001 :  a = '0;
        7'b0011010 :  a = '0;
        7'b0011011 :  a = '0;
        7'b0011100 :  a = '0;
        7'b0011101 :  a = '0;
        7'b0011110 :  a = '0;
        7'b0011111 :  a = '0;
        7'b0100000 :  a = '0;
        7'b0100001 :  a = '0;
        7'b0100010 :  a = '0;
        7'b0100011 :  a = '0;
        7'b0100100 :  a = '0;
        7'b0100101 :  a = '0;
        7'b0100110 :  a = '0;
        7'b0100111 :  a = '0;
        7'b0101000 :  a = '0;
        7'b0101001 :  a = '0;
        7'b0101010 :  a = '0;
        7'b0101011 :  a = '0;
        7'b0101100 :  a = '0;
        7'b0101101 :  a = '0;
        7'b0101110 :  a = '0;
        7'b0101111 :  a = '0;
        7'b0110000 :  a = '0;
        7'b0110001 :  a = '0;
        7'b0110010 :  a = '0;
        7'b0110011 :  a = '0;
        7'b0110100 :  a = '0;
        7'b0110101 :  a = '0;
        7'b0110110 :  a = '0;
        7'b0110111 :  a = '0;
        7'b0111000 :  a = '0;
        7'b0111001 :  a = '0;
        7'b0111010 :  a = '0;
        7'b0111011 :  a = '0;
        7'b0111100 :  a = '0;
        7'b0111101 :  a = '0;
        7'b0111110 :  a = '0;
        7'b0111111 :  a = '0;
        7'b1000000 :  a = '0;
        7'b1000001 :  a = '0;
        7'b1000010 :  a = '0;
        7'b1000011 :  a = '0;
        7'b1000100 :  a = '0;
        7'b1000101 :  a = '0;
        7'b1000110 :  a = '0;
        7'b1000111 :  a = '0;
        7'b1001000 :  a = '0;
        7'b1001001 :  a = '0;
        7'b1001010 :  a = '0;
        7'b1001011 :  a = '0;
        7'b1001100 :  a = '0;
        7'b1001101 :  a = '0;
        7'b1001110 :  a = '0;
        7'b1001111 :  a = '0;
        7'b1010000 :  a = '0;
        7'b1010001 :  a = '0;
        7'b1010010 :  a = '0;
        7'b1010011 :  a = '0;
        7'b1010100 :  a = '0;
        7'b1010101 :  a = '0;
        7'b1010110 :  a = '0;
        7'b1010111 :  a = '0;
        7'b1011000 :  a = '0;
        7'b1011001 :  a = '0;
        7'b1011010 :  a = '0;
        7'b1011011 :  a = '0;
        7'b1011100 :  a = '0;
        7'b1011101 :  a = '0;
        7'b1011110 :  a = '0;
        7'b1011111 :  a = '0;
        7'b1100000 :  a = '0;
        7'b1100001 :  a = '0;
        7'b1100010 :  a = '0;
        7'b1100011 :  a = '0;
        7'b1100100 :  a = '0;
        7'b1100101 :  a = '0;
        7'b1100110 :  a = '0;
        7'b1100111 :  a = '0;
        7'b1101000 :  a = '0;
        7'b1101001 :  a = '0;
        7'b1101010 :  a = '0;
        7'b1101011 :  a = '0;
        7'b1101100 :  a = '0;
        7'b1101101 :  a = '0;
        7'b1101110 :  a = '0;
        7'b1101111 :  a = '0;
        7'b1110000 :  a = '0;
        7'b1110001 :  a = '0;
        7'b1110010 :  a = '0;
        7'b1110011 :  a = '0;
        7'b1110100 :  a = '0;
        7'b1110101 :  a = '0;
        7'b1110110 :  a = '0;
        7'b1110111 :  a = '0;
        7'b1111000 :  a = '0;
        7'b1111001 :  a = '0;
        7'b1111010 :  a = '0;
        7'b1111011 :  a = '0;
        7'b1111100 :  a = '0;
        7'b1111101 :  a = '0;
        7'b1111110 :  a = '0;
        7'b1111111 :  a = '0;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = '0;
        7'b0000001 :  b = '0;
        7'b0000010 :  b = '0;
        7'b0000011 :  b = '0;
        7'b0000100 :  b = '0;
        7'b0000101 :  b = '0;
        7'b0000110 :  b = '0;
        7'b0000111 :  b = '0;
        7'b0001000 :  b = '0;
        7'b0001001 :  b = '0;
        7'b0001010 :  b = '0;
        7'b0001011 :  b = '0;
        7'b0001100 :  b = '0;
        7'b0001101 :  b = '0;
        7'b0001110 :  b = '0;
        7'b0001111 :  b = '0;
        7'b0010000 :  b = '0;
        7'b0010001 :  b = '0;
        7'b0010010 :  b = '0;
        7'b0010011 :  b = '0;
        7'b0010100 :  b = '0;
        7'b0010101 :  b = '0;
        7'b0010110 :  b = '0;
        7'b0010111 :  b = '0;
        7'b0011000 :  b = '0;
        7'b0011001 :  b = '0;
        7'b0011010 :  b = '0;
        7'b0011011 :  b = '0;
        7'b0011100 :  b = '0;
        7'b0011101 :  b = '0;
        7'b0011110 :  b = '0;
        7'b0011111 :  b = '0;
        7'b0100000 :  b = '0;
        7'b0100001 :  b = '0;
        7'b0100010 :  b = '0;
        7'b0100011 :  b = '0;
        7'b0100100 :  b = '0;
        7'b0100101 :  b = '0;
        7'b0100110 :  b = '0;
        7'b0100111 :  b = '0;
        7'b0101000 :  b = '0;
        7'b0101001 :  b = '0;
        7'b0101010 :  b = '0;
        7'b0101011 :  b = '0;
        7'b0101100 :  b = '0;
        7'b0101101 :  b = '0;
        7'b0101110 :  b = '0;
        7'b0101111 :  b = '0;
        7'b0110000 :  b = '0;
        7'b0110001 :  b = '0;
        7'b0110010 :  b = '0;
        7'b0110011 :  b = '0;
        7'b0110100 :  b = '0;
        7'b0110101 :  b = '0;
        7'b0110110 :  b = '0;
        7'b0110111 :  b = '0;
        7'b0111000 :  b = '0;
        7'b0111001 :  b = '0;
        7'b0111010 :  b = '0;
        7'b0111011 :  b = '0;
        7'b0111100 :  b = '0;
        7'b0111101 :  b = '0;
        7'b0111110 :  b = '0;
        7'b0111111 :  b = '0;
        7'b1000000 :  b = '0;
        7'b1000001 :  b = '0;
        7'b1000010 :  b = '0;
        7'b1000011 :  b = '0;
        7'b1000100 :  b = '0;
        7'b1000101 :  b = '0;
        7'b1000110 :  b = '0;
        7'b1000111 :  b = '0;
        7'b1001000 :  b = '0;
        7'b1001001 :  b = '0;
        7'b1001010 :  b = '0;
        7'b1001011 :  b = '0;
        7'b1001100 :  b = '0;
        7'b1001101 :  b = '0;
        7'b1001110 :  b = '0;
        7'b1001111 :  b = '0;
        7'b1010000 :  b = '0;
        7'b1010001 :  b = '0;
        7'b1010010 :  b = '0;
        7'b1010011 :  b = '0;
        7'b1010100 :  b = '0;
        7'b1010101 :  b = '0;
        7'b1010110 :  b = '0;
        7'b1010111 :  b = '0;
        7'b1011000 :  b = '0;
        7'b1011001 :  b = '0;
        7'b1011010 :  b = '0;
        7'b1011011 :  b = '0;
        7'b1011100 :  b = '0;
        7'b1011101 :  b = '0;
        7'b1011110 :  b = '0;
        7'b1011111 :  b = '0;
        7'b1100000 :  b = '0;
        7'b1100001 :  b = '0;
        7'b1100010 :  b = '0;
        7'b1100011 :  b = '0;
        7'b1100100 :  b = '0;
        7'b1100101 :  b = '0;
        7'b1100110 :  b = '0;
        7'b1100111 :  b = '0;
        7'b1101000 :  b = '0;
        7'b1101001 :  b = '0;
        7'b1101010 :  b = '0;
        7'b1101011 :  b = '0;
        7'b1101100 :  b = '0;
        7'b1101101 :  b = '0;
        7'b1101110 :  b = '0;
        7'b1101111 :  b = '0;
        7'b1110000 :  b = '0;
        7'b1110001 :  b = '0;
        7'b1110010 :  b = '0;
        7'b1110011 :  b = '0;
        7'b1110100 :  b = '0;
        7'b1110101 :  b = '0;
        7'b1110110 :  b = '0;
        7'b1110111 :  b = '0;
        7'b1111000 :  b = '0;
        7'b1111001 :  b = '0;
        7'b1111010 :  b = '0;
        7'b1111011 :  b = '0;
        7'b1111100 :  b = '0;
        7'b1111101 :  b = '0;
        7'b1111110 :  b = '0;
        7'b1111111 :  b = '0;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = '0;
        7'b0000001 :  c = '0;
        7'b0000010 :  c = '0;
        7'b0000011 :  c = '0;
        7'b0000100 :  c = '0;
        7'b0000101 :  c = '0;
        7'b0000110 :  c = '0;
        7'b0000111 :  c = '0;
        7'b0001000 :  c = '0;
        7'b0001001 :  c = '0;
        7'b0001010 :  c = '0;
        7'b0001011 :  c = '0;
        7'b0001100 :  c = '0;
        7'b0001101 :  c = '0;
        7'b0001110 :  c = '0;
        7'b0001111 :  c = '0;
        7'b0010000 :  c = '0;
        7'b0010001 :  c = '0;
        7'b0010010 :  c = '0;
        7'b0010011 :  c = '0;
        7'b0010100 :  c = '0;
        7'b0010101 :  c = '0;
        7'b0010110 :  c = '0;
        7'b0010111 :  c = '0;
        7'b0011000 :  c = '0;
        7'b0011001 :  c = '0;
        7'b0011010 :  c = '0;
        7'b0011011 :  c = '0;
        7'b0011100 :  c = '0;
        7'b0011101 :  c = '0;
        7'b0011110 :  c = '0;
        7'b0011111 :  c = '0;
        7'b0100000 :  c = '0;
        7'b0100001 :  c = '0;
        7'b0100010 :  c = '0;
        7'b0100011 :  c = '0;
        7'b0100100 :  c = '0;
        7'b0100101 :  c = '0;
        7'b0100110 :  c = '0;
        7'b0100111 :  c = '0;
        7'b0101000 :  c = '0;
        7'b0101001 :  c = '0;
        7'b0101010 :  c = '0;
        7'b0101011 :  c = '0;
        7'b0101100 :  c = '0;
        7'b0101101 :  c = '0;
        7'b0101110 :  c = '0;
        7'b0101111 :  c = '0;
        7'b0110000 :  c = '0;
        7'b0110001 :  c = '0;
        7'b0110010 :  c = '0;
        7'b0110011 :  c = '0;
        7'b0110100 :  c = '0;
        7'b0110101 :  c = '0;
        7'b0110110 :  c = '0;
        7'b0110111 :  c = '0;
        7'b0111000 :  c = '0;
        7'b0111001 :  c = '0;
        7'b0111010 :  c = '0;
        7'b0111011 :  c = '0;
        7'b0111100 :  c = '0;
        7'b0111101 :  c = '0;
        7'b0111110 :  c = '0;
        7'b0111111 :  c = '0;
        7'b1000000 :  c = '0;
        7'b1000001 :  c = '0;
        7'b1000010 :  c = '0;
        7'b1000011 :  c = '0;
        7'b1000100 :  c = '0;
        7'b1000101 :  c = '0;
        7'b1000110 :  c = '0;
        7'b1000111 :  c = '0;
        7'b1001000 :  c = '0;
        7'b1001001 :  c = '0;
        7'b1001010 :  c = '0;
        7'b1001011 :  c = '0;
        7'b1001100 :  c = '0;
        7'b1001101 :  c = '0;
        7'b1001110 :  c = '0;
        7'b1001111 :  c = '0;
        7'b1010000 :  c = '0;
        7'b1010001 :  c = '0;
        7'b1010010 :  c = '0;
        7'b1010011 :  c = '0;
        7'b1010100 :  c = '0;
        7'b1010101 :  c = '0;
        7'b1010110 :  c = '0;
        7'b1010111 :  c = '0;
        7'b1011000 :  c = '0;
        7'b1011001 :  c = '0;
        7'b1011010 :  c = '0;
        7'b1011011 :  c = '0;
        7'b1011100 :  c = '0;
        7'b1011101 :  c = '0;
        7'b1011110 :  c = '0;
        7'b1011111 :  c = '0;
        7'b1100000 :  c = '0;
        7'b1100001 :  c = '0;
        7'b1100010 :  c = '0;
        7'b1100011 :  c = '0;
        7'b1100100 :  c = '0;
        7'b1100101 :  c = '0;
        7'b1100110 :  c = '0;
        7'b1100111 :  c = '0;
        7'b1101000 :  c = '0;
        7'b1101001 :  c = '0;
        7'b1101010 :  c = '0;
        7'b1101011 :  c = '0;
        7'b1101100 :  c = '0;
        7'b1101101 :  c = '0;
        7'b1101110 :  c = '0;
        7'b1101111 :  c = '0;
        7'b1110000 :  c = '0;
        7'b1110001 :  c = '0;
        7'b1110010 :  c = '0;
        7'b1110011 :  c = '0;
        7'b1110100 :  c = '0;
        7'b1110101 :  c = '0;
        7'b1110110 :  c = '0;
        7'b1110111 :  c = '0;
        7'b1111000 :  c = '0;
        7'b1111001 :  c = '0;
        7'b1111010 :  c = '0;
        7'b1111011 :  c = '0;
        7'b1111100 :  c = '0;
        7'b1111101 :  c = '0;
        7'b1111110 :  c = '0;
        7'b1111111 :  c = '0;
        default    :  c = 'x;
    endcase

	endmodule    
`endif